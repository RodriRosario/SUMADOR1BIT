module C_AND (
  input A,
  input B,
  output OUT
);
  
  assign OUT=A&B;
endmodule